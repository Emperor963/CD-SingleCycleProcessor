module cpu(
    input clk,
    input rst,

    output hlt,
    output [15:0] pc
);


endmodule