module xor (
    input A;
    input B;
    output X;
) ;

assign X = A ^ B;

endmodule