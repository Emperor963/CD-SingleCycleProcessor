module pc_control(
    input B,
    
);

endmodule