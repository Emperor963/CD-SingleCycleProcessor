module paddsb (
    input [15:0] A;
    input [15:0] B;
    input ovfl;

    output []
);

wire [3:0]A_a; //15-12
wire [3:0]A_b; //11-9
wire [3:0]A_c; //8-4
wire [3:0]A_d; //3-0

wire [3:0]B_a; //15-12
wire [3:0]B_b; //11-9
wire [3:0]B_c; //8-4
wire [3:0]B_d; //3-0




assign  = (A_a[3])


endmodule 