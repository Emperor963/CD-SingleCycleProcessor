module ALU(
    input [15:0] In1,
    input [15:0] In2,
    input [2:0] ALUOp,

    output [2:0] FLAG,
    output [15:0] ALUOut
);

wire [15:0] sum;
wire [15:0] difference;
wire [15:0] paddsb;




endmodule