module adder_1bit;

    reg A;
    reg B; 
    reg C;

    wire sum;
    wire overflow;

    




endmodule 