module cpu(
    input clk,
    input rst,

    output hlt,
    output [15:0] pc
);


//Initialize 
wire[2:0] flag_in, flag_out, wr //Flag register variables
wire[15:0] instruction //Instruction wire



endmodule