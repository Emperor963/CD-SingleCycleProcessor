module pc_control(
    input [15:0] pc_in,
    input [8:0] imm,
    input [2:] flags,

    output [15:0] pc_out
);

endmodule